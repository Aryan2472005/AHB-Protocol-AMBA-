module AHB(


          
          );









endmodule
